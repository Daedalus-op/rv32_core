// For slicing the instructions to specific fields
