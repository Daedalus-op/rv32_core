
interface if_id(clk);

endinterface

// --------------------

interface id_eu(clk);

endinterface

// --------------------

interface eu_ma(clk);

endinterface

// --------------------

interface ma_wb(clk);

endinterface
