program rv_test (
	input logic clk
	);
endprogram
