module IF (
    input logic clk,
    input logic 
);
    
endmodule